module Immediate_Generator (
    input  logic [31:0] inst,
    output logic [31:0] imm
);
    // ============================================================
    // Immediate Generator
    // ============================================================
    always_comb begin
        case (inst[6:2])

            // ----------------------------------------------------
            // I-type and Load Instructions
            // ----------------------------------------------------
            `OP_I_LOAD,
            `OP_I_ARITH,
            `OP_JALR,
            `OP_FLW:  imm = {{20{inst[31]}}, inst[31:20]};

            // ----------------------------------------------------
            // S-type and Store Instructions
            // ----------------------------------------------------
            `OP_S_TYPE,
            `OP_FSW:  imm = {{20{inst[31]}}, inst[31:25], inst[11:7]};

            // ----------------------------------------------------
            // B-type
            // ----------------------------------------------------
            `OP_B_TYPE: imm = {{20{inst[31]}}, inst[7], inst[30:25], inst[11:8], 1'b0};

            // ----------------------------------------------------
            // U-type
            // ----------------------------------------------------
            `OP_AUIPC,
            `OP_LUI:  imm = {inst[31:12], 12'd0};

            // ----------------------------------------------------
            // J-type
            // ----------------------------------------------------
            `OP_JAL:  imm = {{12{inst[31]}}, inst[19:12], inst[20],
                             inst[30:25], inst[24:21], 1'b0};

            // ----------------------------------------------------
            // CSR
            // ----------------------------------------------------
            `OP_CSR: imm = {27'd0, inst[19:15]};

            // ----------------------------------------------------
            // Default
            // ----------------------------------------------------
            default:  imm = 32'd0;
        endcase
    end
endmodule
