`include "../include/AXI_define.svh"

module ROM_wrapper (

	input  logic                            clk,
    input  logic                            rst,

    // ReadAddress
    input  logic [`AXI_IDS_BITS-1:0]        ARID_S,
    input  logic [`AXI_ADDR_BITS-1:0]       ARADDR_S,
    input  logic [`AXI_LEN_BITS-1:0]        ARLEN_S,
    input  logic [`AXI_SIZE_BITS-1:0]       ARSIZE_S,
    input  logic [1:0]                      ARBURST_S,
    input  logic                            ARVALID_S,
    output logic                            ARREADY_S,

    // ReadData
    output logic [`AXI_IDS_BITS-1:0]        RID_S,
    output logic [`AXI_DATA_BITS-1:0]       RDATA_S,
    output logic [1:0]                      RRESP_S,
    output logic                            RLAST_S,
    output logic                            RVALID_S,
    input  logic                            RREADY_S,

    // WriteAddress
    input  logic [`AXI_IDS_BITS-1:0]        AWID_S,
    input  logic [`AXI_ADDR_BITS-1:0]       AWADDR_S,
    input  logic [`AXI_LEN_BITS-1:0]        AWLEN_S,
    input  logic [`AXI_SIZE_BITS-1:0]       AWSIZE_S,
    input  logic [1:0]                      AWBURST_S,
    input  logic                            AWVALID_S,
    output logic                            AWREADY_S,

    // WriteData
    input  logic [`AXI_DATA_BITS-1:0]       WDATA_S,
    input  logic [`AXI_STRB_BITS-1:0]       WSTRB_S,
    input  logic                            WLAST_S,
    input  logic                            WVALID_S,
    output logic                            WREADY_S,

    // WriteResponse
    output logic [`AXI_IDS_BITS-1:0]        BID_S,
    output logic [1:0]                      BRESP_S,
    output logic                            BVALID_S,
    input  logic                            BREADY_S,

    // ROM Interface
    output	logic                           ROM_enable,     // CS
    output	logic                           ROM_read,       // OE
    output	logic [11:0]                    ROM_address,    // A
    input	      [`AXI_DATA_BITS-1:0]      ROM_out         // DO
);

	// ============================================================
	// State Definition
	// ============================================================
	typedef enum logic [1:0] {
		ACCEPT        = 2'd0,
		ReadData      = 2'd1,
		WriteData     = 2'd2,
		WriteResponse = 2'd3
	} state_t;

    state_t 				    CurrentState, NextState;

    // ============================================================
	// Local Signals
	// ============================================================
	logic [`AXI_IDS_BITS-1:0] 	AWID, ARID;
	logic [`AXI_DATA_BITS-1:0]  Buffer;
	logic 						Buffer_valid;

	// ============================================================
	// Finite State Machine
	// ============================================================

	// ---------------------------------------
    // State Register
    // ---------------------------------------
	always_ff @( posedge clk or posedge rst ) begin
		if (rst) CurrentState <= ACCEPT;
		else 	 CurrentState <= NextState;
	end

	// ---------------------------------------
    // Next State Logic
    // ---------------------------------------
	always_comb begin
        case(CurrentState)
        ACCEPT: begin
            if      (ARVALID_S) NextState = ReadData;
            else if (AWVALID_S) NextState = WriteData;
            else                NextState = ACCEPT;
        end
        ReadData: begin
            if (RREADY_S)       NextState = ACCEPT;
            else                NextState = CurrentState;
        end
        WriteData: begin
            if (WVALID_S && WLAST_S)
                                NextState = WriteResponse;
            else                NextState = CurrentState;
        end
        WriteResponse: begin
            if(BREADY_S)        NextState = ACCEPT;
            else                NextState = CurrentState;
        end
        endcase
    end

	// ============================================================
    // Channel Output Logic (combinational)
    // ============================================================
    always_comb begin
        ARREADY_S = 1'b0;
        AWREADY_S = 1'b0;
        RID_S     = `AXI_IDS_BITS'd0;
        RDATA_S   = `AXI_DATA_BITS'd0;
        RRESP_S   = `AXI_RESP_DECERR;
        RVALID_S  = 1'b0;
        RLAST_S   = 1'b0;
        WREADY_S  = 1'b0;
        BID_S     = `AXI_IDS_BITS'd0;
        BVALID_S  = 1'b0;
        BRESP_S   = `AXI_RESP_DECERR;

        case (CurrentState)
            ACCEPT: begin
                ARREADY_S = 1'b1;
                AWREADY_S = 1'b1;
            end
            ReadData: begin
                RID_S     = ARID;
                RDATA_S   = (Buffer_valid) ? Buffer : ROM_out;
                RRESP_S   = `AXI_RESP_OKAY;
                RVALID_S  = 1'b1;
                RLAST_S   = 1'b1;
            end
            WriteData: begin
                WREADY_S  = 1'b1;
            end
            WriteResponse: begin
                BID_S     = AWID;
                BVALID_S  = 1'b1;
                BRESP_S   = `AXI_RESP_SLVERR;
            end
        endcase
    end

	// ============================================================
	// ID Storage
	// ============================================================
	always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            ARID  <= `AXI_IDS_BITS'd0;
            AWID  <= `AXI_IDS_BITS'd0;
        end
        else if (CurrentState == ACCEPT) begin
            ARID  <= ARVALID_S ? ARID_S : ARID;
            AWID  <= AWVALID_S ? AWID_S : AWID;
        end
    end

    // ============================================================
	// Read Data Buffer
	// ============================================================
	always_ff @( posedge clk or posedge rst ) begin // Waiting
		if (rst) begin
            Buffer_valid <= 1'b0;
            Buffer       <= `AXI_DATA_BITS'd0;
        end else if (CurrentState == ReadData) begin
            if (RREADY_S && RVALID_S) begin
                Buffer_valid <= 1'b0;
                Buffer       <= `AXI_DATA_BITS'd0;
            end else begin
                Buffer_valid <= 1'b1;
                Buffer       <= ROM_out;
            end
		end
	end

    // ============================================================
	// ROM Interface
	// ============================================================
    always_comb begin
        case (CurrentState)
            ACCEPT : begin
                ROM_enable  = ARVALID_S;
                ROM_read    = 1'b0;
                ROM_address = ARVALID_S ? ARADDR_S[13:2] : 12'd0;
            end
            ReadData : begin
                ROM_enable  = 1'b0;
                ROM_read    = 1'b1;
                ROM_address = 12'd0;
            end
            default : begin
                ROM_enable  = 1'b0;
                ROM_read    = 1'b0;
                ROM_address = 12'd0;
            end
        endcase
    end



endmodule